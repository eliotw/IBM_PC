
module 75477(
	     a,
	     y
	     );

   input [1:0] a;
   output [1:0] y;

endmodule // 75477
