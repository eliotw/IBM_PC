
module ls245(
	     a,
	     b,
	     dir,
	     g_n
	     );

   inout [7:0] a;
   inout [7:0] b;
   input       dir;
   input       g_n;

endmodule // ls245
