
module ls158(
	     a,
	     b,
	     y,
	     s,
	     g
	     );

   input [3:0] a, b;
   input       s, g;
   output [3:0] y;

endmodule // ls158
