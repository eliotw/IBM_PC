
module ls244(
	     a,
	     y,
	     g1_n,
	     g2_n);

   inout [7:0] a;
   inout [7:0] y;
   input       g1_n, g2_n;

endmodule // ls244
