/*
 * sdcard:
 * Verilog description of module that mimics the SD card reader in the ao486
 * floppy disk file
 */

module sdcard(
	      // inputs go here
	      );

   // Wires

   // Registers

   // Assignments

   // Block RAM

endmodule // sdcard
