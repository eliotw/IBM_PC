
module ls322(
	     q,
	     qh1,
	     oe_n,
	     di,
	     do,
	     clr_n,
	     clock,
	     se_n,
	     ds,
	     sp_n,
	     g_n
	     );

   input [7:0] q;
   output      qh1;
   input       oe_n, di, do, clr_n, clock, se_n, ds, sp_n, g_n;

endmodule // ls322
