
module rds(
	   // ?
	   );

endmodule // rds
