
module ls670(
	     d,
	     q,
	     ra,
	     rb,
	     read,
	     wa,
	     wb,
	     write
	     );

   input [3:0] d;
   output [3:0] q;
   input 	ra, rb, read, wa, wb, write;

endmodule // ls670
