library verilog;
use verilog.vl_types.all;
entity test_zet is
end test_zet;
