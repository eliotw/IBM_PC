
module ls138(
	     a, b, c,
	     g2b, g2a,
	     g1,
	     y
	     );

   output [7:0] y;
   input 	a, b, c, g2b, g2a, g1;

endmodule // ls138
