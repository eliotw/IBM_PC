
module timedelay(
		 in,
		 t25,
		 t75,
		 t125
		 );

   input in;
   output t25, t75, t125;

endmodule // timedelay
