// PLEASE SEE MODULE LS280 UNDER "RAM" FOLDER

module s280(
	    md,
	    i,
	    odd,
	    even
	    );

   input [7:0] md;
   input       i;
   output      odd, even;

endmodule // s280
