// MOVED TO RAM FOLDER
module rds(
	   // ?
	   );

endmodule // rds
