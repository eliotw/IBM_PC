
module ls373(
	     d,
	     q,
	     g,
	     oe_n
	     );

   inout [7:0] d;
   inout [7:0] q;
   input       g;
   input       oe_n;

endmodule // ls373
